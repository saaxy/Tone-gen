library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Tone_Generator is
    Port (
        clk : in STD_LOGIC;
        en : in STD_LOGIC;
        tone_freq : in STD_LOGIC_VECTOR (4 downto 0);
        tone_ampl : in STD_LOGIC_VECTOR (3 downto 0); -- change by 1/15 of volume
        pwm_out : out STD_LOGIC
    );
end Tone_Generator;

architecture Behavioral of Tone_Generator is
    signal counter : integer := 1;
    signal threshold : integer := 1;
   
    signal i : integer :=1;
    signal decoded_points : integer := 0;
   
    type Frequency_array is array (1 to 32) of integer;
    signal F_Array : Frequency_array := (2616, 2937, 3296, 3492, 3920, 4400, 4939, 5233, 5873, 6593, 6985, 7840, 8800, 9878, 10470, 11750, 13190,13970 , 15680, 17600, 19760, 20930, 23490, 26370, 27940, 31360, 35200, 39510, 41860, 46990, 52740, 55880); -- 10x bigger than original, to not use float C2 -> G4
       

    signal Amplitude : integer := 1;
   
   
    constant zero : integer := 500;
    constant divided_points : integer := 1024 ;
    type Time_array is array(1 to divided_points) of Integer;
    signal T_array : Time_array := (0,3,6,9,12,15,18,21,25,28,31,34,37,40,43,46,49,52,55,58,61,64,67,70,73,76,79,82,85,89,92,95,98,101,104,107,110,113,116,119,121,124,127,130,133,136,139,142,145,148,151,154,157,160,163,166,168,171,174,177,180,183,186,189,191,194,197,200,203,205,208,211,214,217,219,222,225,228,230,233,236,238,241,244,246,249,252,254,257,260,262,265,267,270,273,275,278,280,283,285,288,290,293,295,298,300,303,305,308,310,312,315,317,320,322,324,327,329,331,333,336,338,340,343,345,347,349,351,354,356,358,360,362,364,366,368,370,373,375,377,379,381,383,385,387,388,390,392,394,396,398,400,402,403,405,407,409,411,412,414,416,417,419,421,422,424,426,427,429,430,432,434,435,437,438,440,441,442,444,445,447,448,449,451,452,453,455,456,457,458,460,461,462,463,464,465,466,468,469,470,471,472,473,474,475,476,477,478,478,479,480,481,482,483,483,484,485,486,486,487,488,489,489,490,490,491,492,492,493,493,494,494,495,495,495,496,496,497,497,497,498,498,498,498,499,499,499,499,499,500,500,500,500,500,500,500,500,500,500,500,500,500,500,500,499,499,499,499,499,498,498,498,498,497,497,497,496,496,495,495,495,494,494,493,493,492,492,491,490,490,489,489,488,487,486,486,485,484,483,483,482,481,480,479,478,478,477,476,475,474,473,472,471,470,469,468,466,465,464,463,462,461,460,458,457,456,455,453,452,451,449,448,447,445,444,442,441,440,438,437,435,434,432,430,429,427,426,424,422,421,419,417,416,414,412,411,409,407,405,403,402,400,398,396,394,392,390,388,387,385,383,381,379,377,375,373,370,368,366,364,362,360,358,356,354,351,349,347,345,343,340,338,336,333,331,329,327,324,322,320,317,315,312,310,308,305,303,300,298,295,293,290,288,285,283,280,278,275,273,270,267,265,262,260,257,254,252,249,246,244,241,238,236,233,230,228,225,222,219,217,214,211,208,205,203,200,197,194,191,189,186,183,180,177,174,171,168,166,163,160,157,154,151,148,145,142,139,136,133,130,127,124,121,119,116,113,110,107,104,101,98,95,92,89,85,82,79,76,73,70,67,64,61,58,55,52,49,46,43,40,37,34,31,28,25,21,18,15,12,9,6,3,0,-3,-6,-9,-12,-15,-18,-21,-25,-28,-31,-34,-37,-40,-43,-46,-49,-52,-55,-58,-61,-64,-67,-70,-73,-76,-79,-82,-85,-89,-92,-95,-98,-101,-104,-107,-110,-113,-116,-119,-121,-124,-127,-130,-133,-136,-139,-142,-145,-148,-151,-154,-157,-160,-163,-166,-168,-171,-174,-177,-180,-183,-186,-189,-191,-194,-197,-200,-203,-205,-208,-211,-214,-217,-219,-222,-225,-228,-230,-233,-236,-238,-241,-244,-246,-249,-252,-254,-257,-260,-262,-265,-267,-270,-273,-275,-278,-280,-283,-285,-288,-290,-293,-295,-298,-300,-303,-305,-308,-310,-312,-315,-317,-320,-322,-324,-327,-329,-331,-333,-336,-338,-340,-343,-345,-347,-349,-351,-354,-356,-358,-360,-362,-364,-366,-368,-370,-373,-375,-377,-379,-381,-383,-385,-387,-388,-390,-392,-394,-396,-398,-400,-402,-403,-405,-407,-409,-411,-412,-414,-416,-417,-419,-421,-422,-424,-426,-427,-429,-430,-432,-434,-435,-437,-438,-440,-441,-442,-444,-445,-447,-448,-449,-451,-452,-453,-455,-456,-457,-458,-460,-461,-462,-463,-464,-465,-466,-468,-469,-470,-471,-472,-473,-474,-475,-476,-477,-478,-478,-479,-480,-481,-482,-483,-483,-484,-485,-486,-486,-487,-488,-489,-489,-490,-490,-491,-492,-492,-493,-493,-494,-494,-495,-495,-495,-496,-496,-497,-497,-497,-498,-498,-498,-498,-499,-499,-499,-499,-499,-500,-500,-500,-500,-500,-500,-500,-500,-500,-500,-500,-500,-500,-500,-500,-499,-499,-499,-499,-499,-498,-498,-498,-498,-497,-497,-497,-496,-496,-495,-495,-495,-494,-494,-493,-493,-492,-492,-491,-490,-490,-489,-489,-488,-487,-486,-486,-485,-484,-483,-483,-482,-481,-480,-479,-478,-478,-477,-476,-475,-474,-473,-472,-471,-470,-469,-468,-466,-465,-464,-463,-462,-461,-460,-458,-457,-456,-455,-453,-452,-451,-449,-448,-447,-445,-444,-442,-441,-440,-438,-437,-435,-434,-432,-430,-429,-427,-426,-424,-422,-421,-419,-417,-416,-414,-412,-411,-409,-407,-405,-403,-402,-400,-398,-396,-394,-392,-390,-388,-387,-385,-383,-381,-379,-377,-375,-373,-370,-368,-366,-364,-362,-360,-358,-356,-354,-351,-349,-347,-345,-343,-340,-338,-336,-333,-331,-329,-327,-324,-322,-320,-317,-315,-312,-310,-308,-305,-303,-300,-298,-295,-293,-290,-288,-285,-283,-280,-278,-275,-273,-270,-267,-265,-262,-260,-257,-254,-252,-249,-246,-244,-241,-238,-236,-233,-230,-228,-225,-222,-219,-217,-214,-211,-208,-205,-203,-200,-197,-194,-191,-189,-186,-183,-180,-177,-174,-171,-168,-166,-163,-160,-157,-154,-151,-148,-145,-142,-139,-136,-133,-130,-127,-124,-121,-119,-116,-113,-110,-107,-104,-101,-98,-95,-92,-89,-85,-82,-79,-76,-73,-70,-67,-64,-61,-58,-55,-52,-49,-46,-43,-40,-37,-34,-31,-28,-25,-21,-18,-15,-12,-9,-6,-3);
    
    begin

      freq_decoder: process (tone_freq) -- decoding frequencies
    begin
        case tone_freq is
            when "00000" =>    
                decoded_points <= 1_000_000_000 / (F_array(1)*divided_points);
            when "00001" =>    
                decoded_points <= 1000000000 / (F_array(2)*divided_points);
            when "00010" =>    
                decoded_points <= 1000000000 / (F_array(3)*divided_points);
            when "00011" =>    
                decoded_points <= 1000000000 / (F_array(4)*divided_points);
            when "00100" =>    
                decoded_points <= 1000000000 / (F_array(5)*divided_points);
            when "00101" =>    
                decoded_points <= 1000000000 / (F_array(6)*divided_points);
            when "00110" =>    
                decoded_points <= 1000000000 / (F_array(7)*divided_points);  
            when "00111" =>    
                decoded_points <= 1000000000 / (F_array(8)*divided_points);  
            when "01000" =>    
                decoded_points <= 1000000000 / (F_array(9)*divided_points);
            when "01001" =>    
                decoded_points <= 1000000000 / (F_array(10)*divided_points);
            when "01010" =>    
                decoded_points <= 1000000000 / (F_array(11)*divided_points);
            when "01011" =>    
                decoded_points <= 1000000000 / (F_array(12)*divided_points);
            when "01100" =>    
                decoded_points <= 1000000000 / (F_array(13)*divided_points);
            when "01101" =>    
                decoded_points <= 1000000000 / (F_array(14)*divided_points);
            when "01110" =>    
                decoded_points <= 1000000000 / (F_array(15)*divided_points);
            when "01111" =>    
                decoded_points <= 1000000000 / (F_array(16)*divided_points);
            when "10000" =>    
                decoded_points <= 1000000000 / (F_array(17)*divided_points);  
            when "10001" =>    
                decoded_points <= 1000000000 / (F_array(18)*divided_points);  
            when "10010" =>    
                decoded_points <= 1000000000 / (F_array(19)*divided_points);
            when "10011" =>    
                decoded_points <= 1000000000 / (F_array(20)*divided_points);
            when "10100" =>    
                decoded_points <= 1000000000 / (F_array(21)*divided_points);
            when "10101" =>    
                decoded_points <= 1000000000 / (F_array(22)*divided_points);
            when "10110" =>    
                decoded_points <= 1000000000 / (F_array(23)*divided_points);
            when "10111" =>    
                decoded_points <= 1000000000 / (F_array(24)*divided_points);
            when "11000" =>    
                decoded_points <= 1000000000 / (F_array(25)*divided_points);
            when "11001" =>    
                decoded_points <= 1000000000 / (F_array(26)*divided_points);
            when "11010" =>    
                decoded_points <= 1000000000 / (F_array(27)*divided_points);  
            when "11011" =>    
                decoded_points <= 1000000000 / (F_array(28)*divided_points);  
            when "11100" =>    
                decoded_points <= 1000000000 / (F_array(29)*divided_points);
            when "11101" =>    
                decoded_points <= 1000000000 / (F_array(30)*divided_points);
            when "11110" =>    
                decoded_points <= 1000000000 / (F_array(31)*divided_points);
            when "11111" =>    
                decoded_points <= 1000000000 / (F_array(32)*divided_points);
            when others =>
                decoded_points <= 0;
        end case;
    end process;
   
    amplitude_decoder: process (tone_ampl) -- decoding amplitude
    begin
        Amplitude <= (1000 * to_integer(unsigned(tone_ampl))) / 15;
    end process;
   
    process (clk, en, i) -- generating PWM to sinewave
    begin
        if en = '0' then
            counter <= 0;
            pwm_out <= '0';
        else
            threshold <= (((T_array(i) * Amplitude)/1000 + zero) * decoded_points/1000);
            if rising_edge(clk) then
                  counter <= counter + 1;
                if counter >= decoded_points then
                    i <= i + 1;
                    if i >= divided_points then
                    i <= 1;
                    end if;
                    counter <= 0;
                end if;
                if counter < threshold then
                  pwm_out <= '1';
                  else
                  pwm_out <= '0';
                  end if;
            end if;
        end if;
    end process;
   
end Behavioral;